// ------------------------------------------------------------------------------------------------
// Copyright 2022 by Heqing Huang (feipenghhq@gamil.com)
// Author: Heqing Huang
//
// Date Created: 01/17/2022
// ------------------------------------------------------------------------------------------------
// veriRISCV
// ------------------------------------------------------------------------------------------------
// Define file for veriRISCV core
// ------------------------------------------------------------------------------------------------


`ifndef _VERIRISCV_CORE_
`define _VERIRISCV_CORE_


`include "core_arch.svh"
`include "core_struct.svh"
`include "core_opcode.svh"

`endif
